`define MODULE_NAME Square_linear_div
`define UNSIGNED
`define NO_REMAINDER
