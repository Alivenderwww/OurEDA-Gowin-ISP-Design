parameter M=34;
parameter N=42;
parameter LATENCY=20;
