`define MODULE_NAME Hue_Cal_Division
`define UNSIGNED
`define NO_REMAINDER
