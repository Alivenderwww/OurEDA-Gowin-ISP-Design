`define MODULE_NAME AWB_Integer_Division
`define UNSIGNED
`define NO_REMAINDER
