`define MODULE_NAME Sat_Cal_Division
`define UNSIGNED
`define NO_REMAINDER
