parameter M=8;
parameter N=16;
parameter LATENCY=5;
