parameter M=11;
parameter N=17;
parameter LATENCY=5;
